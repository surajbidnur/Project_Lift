library verilog;
use verilog.vl_types.all;
entity liftsm_tb is
end liftsm_tb;
